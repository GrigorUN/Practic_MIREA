library verilog;
use verilog.vl_types.all;
entity LAB_3_vlg_vec_tst is
end LAB_3_vlg_vec_tst;
