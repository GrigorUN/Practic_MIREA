library verilog;
use verilog.vl_types.all;
entity LAB_4_2_vlg_vec_tst is
end LAB_4_2_vlg_vec_tst;
