library verilog;
use verilog.vl_types.all;
entity LAB_2_1 is
    port(
        LESS            : out    vl_logic;
        B1              : in     vl_logic;
        A1              : in     vl_logic;
        B2              : in     vl_logic;
        A2              : in     vl_logic;
        B0              : in     vl_logic;
        A0              : in     vl_logic
    );
end LAB_2_1;
