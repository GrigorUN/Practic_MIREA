library verilog;
use verilog.vl_types.all;
entity LAB1_1_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LAB1_1_vlg_check_tst;
