library verilog;
use verilog.vl_types.all;
entity LAB_1_2_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LAB_1_2_vlg_check_tst;
