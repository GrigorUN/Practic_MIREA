library verilog;
use verilog.vl_types.all;
entity LAB_3_vlg_check_tst is
    port(
        LESS            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LAB_3_vlg_check_tst;
