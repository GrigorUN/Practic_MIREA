library verilog;
use verilog.vl_types.all;
entity LAB_2_1_vlg_vec_tst is
end LAB_2_1_vlg_vec_tst;
