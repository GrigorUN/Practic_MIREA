library verilog;
use verilog.vl_types.all;
entity LAB1_1 is
    port(
        Y               : out    vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic
    );
end LAB1_1;
