library verilog;
use verilog.vl_types.all;
entity LAB_2_2 is
    port(
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        b0              : in     vl_logic;
        b1              : in     vl_logic;
        b2              : in     vl_logic;
        y               : out    vl_logic
    );
end LAB_2_2;
