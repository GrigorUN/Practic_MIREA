library verilog;
use verilog.vl_types.all;
entity LAB1_1_vlg_vec_tst is
end LAB1_1_vlg_vec_tst;
